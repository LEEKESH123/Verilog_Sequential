module SR_ff(rst,clk,s,r,q,qbar);
	input rst,clk,s,r;
	output reg q;
	output qbar;
	assign qbar = ~q;
	always@(posedge clk or posedge rst) begin
	if(rst)
		q <= 0;
	else begin
		case ({s,r})
		2'b00 : q <= q;
		2'b01 : q <= 0;
		2'b10 : q <= 1;
		default : q=1'bZ;
		endcase
		end
	end
endmodule
